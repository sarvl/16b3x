LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY ram IS
	PORT(
		a0  : IN  std_logic_vector(15 DOWNTO 0);
		i0  : IN  std_logic_vector(15 DOWNTO 0);
		o0  : OUT std_logic_vector(15 DOWNTO 0);

		we  : IN  std_logic := '0';
		clk : IN  std_logic);
END ENTITY ram;

ARCHITECTURE behav OF RAM IS 
	TYPE arr IS ARRAY(32767 DOWNTO 0) OF std_logic_vector(7 DOWNTO 0);
	SIGNAL datam : arr := (
	--fib.asm
	-- 00 => x"28", 01 => x"29", 02 => x"2F", 03 => x"8F", 04 => x"A6", 
	-- 05 => x"02", 06 => x"00", 07 => x"01", 08 => x"CF", 09 => x"A3", 
	-- 10 => x"38", 11 => x"00", 12 => x"0F",
	--fact.asm
	-- 00 => x"A7", 01 => x"89", 02 => x"A5", 03 => x"28", 04 => x"A7", 
	-- 05 => x"02", 06 => x"C9", 07 => x"00", 08 => x"C9", 09 => x"A1", 
	-- 10 => x"B7", 11 => x"07", 12 => x"77", 13 => x"88", 14 => x"A6", 
	-- 15 => x"70", 16 => x"C8", 17 => x"AB", 18 => x"79", 19 => x"AF", 
	-- 20 => x"A7", 21 => x"28", 22 => x"7F", 23 => x"02", 24 => x"B7", 
	-- 25 => x"28", 26 => x"AF", 27 => x"38", 28 => x"0F",
	--sort.asm
	00 => x"A7", 01 => x"89", 02 => x"A5", 03 => x"28", 04 => x"A7", 
	05 => x"02", 06 => x"C9", 07 => x"00", 08 => x"C9", 09 => x"A1", 
	10 => x"B7", 11 => x"8A", 12 => x"B6", 13 => x"03", 14 => x"03", 
	15 => x"C0", 16 => x"C1", 17 => x"CA", 18 => x"A7", 19 => x"06", 
	20 => x"06", 21 => x"89", 22 => x"B6", 23 => x"02", 24 => x"03", 
	25 => x"C3", 26 => x"04", 27 => x"05", 28 => x"04", 29 => x"A6", 
	30 => x"05", 31 => x"04", 32 => x"C2", 33 => x"C3", 34 => x"03",
	35 => x"A4", 36 => x"C9", 37 => x"A1", 38 => x"B7", 39 => x"2E",
	40 => x"28", 41 => x"29", 42 => x"AF", 43 => x"F0", 44 => x"F8", 
	45 => x"00", 46 => x"CE", 47 => x"8E", 48 => x"A3", 49 => x"28", 
	50 => x"29", 51 => x"2A", 52 => x"AF", 53 => x"28", 54 => x"29", 
	55 => x"AF", 56 => x"30", 57 => x"31", 58 => x"32", 59 => x"33", 
	60 => x"34", 61 => x"35", 62 => x"36", 63 => x"37", 64 => x"0F",
	--pipeline_easy.asm
	-- 00 => x"28", 01 => x"29", 02 => x"2A", 03 => x"2B", 04 => x"2C", 
	-- 05 => x"2D", 06 => x"2E", 07 => x"2F", 08 => x"00", 09 => x"01", 
	-- 10 => x"02", 11 => x"03", 12 => x"04", 13 => x"05", 14 => x"06", 
	-- 15 => x"07", 16 => x"F0", 17 => x"F1", 18 => x"F2", 19 => x"F3", 
	-- 20 => x"F4", 21 => x"F5", 22 => x"F6", 23 => x"F7", 24 => x"0F",
	--pipeline_alu_dep.asm
	-- 00 => x"29", 01 => x"28", 02 => x"F0", 03 => x"02", 04 => x"F8",
	-- 05 => x"03", 06 => x"C0", 07 => x"C8", 08 => x"F8", 09 => x"04",
	-- 10 => x"0F",

		OTHERS => x"00"
	);
	SIGNAL datal : arr := (
	--fib.asm
	-- 00 => x"00", 01 => x"01", 02 => x"07", 03 => x"00", 04 => x"0A", 
	-- 05 => x"05", 06 => x"25", 07 => x"58", 08 => x"01", 09 => x"05", 
	-- 10 => x"50", 11 => x"00", 12 => x"00", 
	--fact.asm
	-- 00 => x"19", 01 => x"00", 02 => x"05", 03 => x"00", 04 => x"0A", 
	-- 05 => x"05", 06 => x"01", 07 => x"58", 08 => x"01", 09 => x"07", 
	-- 10 => x"00", 11 => x"4C", 12 => x"00", 13 => x"01", 14 => x"15", 
	-- 15 => x"00", 16 => x"01", 17 => x"0B", 18 => x"00", 19 => x"01", 
	-- 20 => x"16", 21 => x"01", 22 => x"00", 23 => x"ED", 24 => x"00", 
	-- 25 => x"06", 26 => x"0B", 27 => x"50", 28 => x"00",
	--sort.asm
	00 => x"27", 01 => x"00", 02 => x"05", 03 => x"00", 04 => x"0A", 
	05 => x"05", 06 => x"01", 07 => x"58", 08 => x"01", 09 => x"07", 
	10 => x"00", 11 => x"00", 12 => x"00", 13 => x"06", 14 => x"27", 
	15 => x"02", 16 => x"02", 17 => x"02", 18 => x"0B", 19 => x"05", 
	20 => x"38", 21 => x"02", 22 => x"00", 23 => x"05", 24 => x"05", 
	25 => x"02", 26 => x"46", 27 => x"66", 28 => x"B1", 29 => x"20", 
	30 => x"47", 31 => x"67", 32 => x"02", 33 => x"02", 34 => x"D1",
	35 => x"1A", 36 => x"02", 37 => x"13", 38 => x"00", 39 => x"A4", 
	40 => x"01", 41 => x"7B", 42 => x"01", 43 => x"01", 44 => x"01", 
	45 => x"C7", 46 => x"02", 47 => x"96", 48 => x"29", 49 => x"96", 
	50 => x"C8", 51 => x"10", 52 => x"0B", 53 => x"96", 54 => x"10", 
	55 => x"13", 56 => x"96", 57 => x"98", 58 => x"9A", 59 => x"9C", 
	60 => x"9E", 61 => x"A0", 62 => x"A2", 63 => x"A4", 64 => x"00",
	--pipeline_easy.asm
	-- 00 => x"00", 01 => x"01", 02 => x"02", 03 => x"03", 04 => x"04", 
	-- 05 => x"05", 06 => x"06", 07 => x"07", 08 => x"38", 09 => x"58", 
	-- 10 => x"78", 11 => x"98", 12 => x"B8", 13 => x"D8", 14 => x"F8", 
	-- 15 => x"18", 16 => x"01", 17 => x"01", 18 => x"01", 19 => x"01", 
	-- 20 => x"01", 21 => x"01", 22 => x"01", 23 => x"01", 24 => x"00",
	--pipeline_alu_dep.asm
	-- 00 => x"00", 01 => x"10", 02 => x"02", 03 => x"05", 04 => x"02",
	-- 05 => x"05", 06 => x"01", 07 => x"02", 08 => x"01", 09 => x"05",
	-- 10 => x"00",
		
		OTHERS => x"00"
	);

	SIGNAL a0m : std_logic_vector(14 DOWNTO 0);
	SIGNAL a0l : std_logic_vector(14 DOWNTO 0);
	
BEGIN
	a0m <= a0(15 DOWNTO 1);
	a0l <= a0(15 DOWNTO 1);

	datam(to_integer(unsigned(a0m))) <= i0(15 DOWNTO 8) WHEN we = '1' AND rising_edge(clk);
	datal(to_integer(unsigned(a0l))) <= i0( 7 DOWNTO 0) WHEN we = '1' AND rising_edge(clk);

	o0 <= datam(to_integer(unsigned(a0m))) 
	    & datal(to_integer(unsigned(a0l)));


END ARCHITECTURE behav;
